-- tug.vhd: Module to implement a game of Tug of War in VHDL
-- todo: finish this
