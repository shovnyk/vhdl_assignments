-- magcomp_tb.vhd: Testbench to test a 4 bit magnitude comparator


