-- counter_control_tb.vhd: Testbench to test the counter module
-- todo: finish this

library ieee;
use ieee.std_logic_1164.all;

entity counter_control_tb is
end counter_control_tb;

architecture sim of counter_control_tb is
begin
end sim;
