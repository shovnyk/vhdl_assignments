-- park_tb.vhd: Test bench to test the car parking FSM
-- todo : finish this

library ieee;
use ieee.std_logic_1164.all;
