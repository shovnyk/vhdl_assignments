-- fsm15_tb.vhd: Testbench to test the FSM in question 15
-- todo finish this
