-- fsm16_tb.vhd: Testbench to test the FSM in question 16
-- todo: finish this
