-- debounce.vhd: Module to debounce a push buttong switch
-- todo: finish this

entity debouncer is 
end debouncer;

architecture behavioral of debouncer is
begin
end behavioral;
